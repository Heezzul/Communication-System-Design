library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;


package mypackage is
   type std_2b_array is array(natural range <>) of std_logic_vector(1 downto 0);
   type std_3b_array is array(natural range <>) of std_logic_vector(2 downto 0);
   type std_4b_array is array(natural range <>) of std_logic_vector(3 downto 0);
   type std_5b_array is array(natural range <>) of std_logic_vector(4 downto 0);
   type std_6b_array is array(natural range <>) of std_logic_vector(5 downto 0);
   type std_7b_array is array(natural range <>) of std_logic_vector(6 downto 0);
   type std_8b_array is array(natural range <>) of std_logic_vector(7 downto 0);
   type std_9b_array is array(natural range <>) of std_logic_vector(8 downto 0);
   type std_10b_array is array(natural range <>) of std_logic_vector(9 downto 0);
   type std_11b_array is array(natural range <>) of std_logic_vector(10 downto 0);
   type std_12b_array is array(natural range <>) of std_logic_vector(11 downto 0);
   type std_13b_array is array(natural range <>) of std_logic_vector(12 downto 0);
   type std_14b_array is array(natural range <>) of std_logic_vector(13 downto 0);
   type std_15b_array is array(natural range <>) of std_logic_vector(14 downto 0);
   type std_16b_array is array(natural range <>) of std_logic_vector(15 downto 0);
   type std_17b_array is array(natural range <>) of std_logic_vector(16 downto 0);
   type std_18b_array is array(natural range <>) of std_logic_vector(17 downto 0);
   type std_19b_array is array(natural range <>) of std_logic_vector(18 downto 0);
   type std_20b_array is array(natural range <>) of std_logic_vector(19 downto 0);
   type std_21b_array is array(natural range <>) of std_logic_vector(20 downto 0);
   type std_22b_array is array(natural range <>) of std_logic_vector(21 downto 0);
   type std_23b_array is array(natural range <>) of std_logic_vector(22 downto 0);
   type std_24b_array is array(natural range <>) of std_logic_vector(23 downto 0);
   type std_25b_array is array(natural range <>) of std_logic_vector(24 downto 0);  
end mypackage;


package body mypackage is
end mypackage;

