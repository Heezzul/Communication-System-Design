library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;

package NCO_ROM_package is
		constant NCOROM_Address : integer := 2**8;
		constant NCOROM_Data : integer := 10;
		
		Type ROM_TYPE is array(0 to 255) of std_logic_vector(9 downto 0);
		
		constant COSROM_Table : ROM_TYPE := ROM_TYPE '( 		

  				conv_std_logic_vector( 511 , 10),
  				conv_std_logic_vector( 511 , 10),
  				conv_std_logic_vector( 510 , 10),
  				conv_std_logic_vector( 510 , 10),
  				conv_std_logic_vector( 509 , 10),
  				conv_std_logic_vector( 507 , 10),
  				conv_std_logic_vector( 505 , 10),
  				conv_std_logic_vector( 503 , 10),
  				conv_std_logic_vector( 501 , 10),
  				conv_std_logic_vector( 499 , 10),
  				conv_std_logic_vector( 496 , 10),
  				conv_std_logic_vector( 492 , 10),
  				conv_std_logic_vector( 489 , 10),
  				conv_std_logic_vector( 485 , 10),
  				conv_std_logic_vector( 481 , 10),
  				conv_std_logic_vector( 477 , 10),
  				conv_std_logic_vector( 472 , 10),
  				conv_std_logic_vector( 467 , 10),
  				conv_std_logic_vector( 462 , 10),
  				conv_std_logic_vector( 456 , 10),
  				conv_std_logic_vector( 451 , 10),
  				conv_std_logic_vector( 445 , 10),
  				conv_std_logic_vector( 438 , 10),
  				conv_std_logic_vector( 432 , 10),
  				conv_std_logic_vector( 425 , 10),
  				conv_std_logic_vector( 418 , 10),
  				conv_std_logic_vector( 410 , 10),
  				conv_std_logic_vector( 403 , 10),
  				conv_std_logic_vector( 395 , 10),
  				conv_std_logic_vector( 387 , 10),
  				conv_std_logic_vector( 379 , 10),
  				conv_std_logic_vector( 370 , 10),
  				conv_std_logic_vector( 361 , 10),
  				conv_std_logic_vector( 352 , 10),
  				conv_std_logic_vector( 343 , 10),
  				conv_std_logic_vector( 334 , 10),
  				conv_std_logic_vector( 324 , 10),
  				conv_std_logic_vector( 314 , 10),
  				conv_std_logic_vector( 304 , 10),
  				conv_std_logic_vector( 294 , 10),
  				conv_std_logic_vector( 284 , 10),
  				conv_std_logic_vector( 273 , 10),
  				conv_std_logic_vector( 263 , 10),
  				conv_std_logic_vector( 252 , 10),
  				conv_std_logic_vector( 241 , 10),
  				conv_std_logic_vector( 230 , 10),
  				conv_std_logic_vector( 218 , 10),
  				conv_std_logic_vector( 207 , 10),
  				conv_std_logic_vector( 196 , 10),
  				conv_std_logic_vector( 184 , 10),
  				conv_std_logic_vector( 172 , 10),
  				conv_std_logic_vector( 160 , 10),
  				conv_std_logic_vector( 148 , 10),
  				conv_std_logic_vector( 136 , 10),
  				conv_std_logic_vector( 124 , 10),
  				conv_std_logic_vector( 112 , 10),
  				conv_std_logic_vector( 100 , 10),
  				conv_std_logic_vector(  87 , 10),
  				conv_std_logic_vector(  75 , 10),
  				conv_std_logic_vector(  63 , 10),
  				conv_std_logic_vector(  50 , 10),
  				conv_std_logic_vector(  38 , 10),
  				conv_std_logic_vector(  25 , 10),
  				conv_std_logic_vector(  13 , 10),
  				conv_std_logic_vector(   0 , 10),
  				conv_std_logic_vector( -13 , 10),
  				conv_std_logic_vector( -25 , 10),
  				conv_std_logic_vector( -38 , 10),
  				conv_std_logic_vector( -50 , 10),
  				conv_std_logic_vector( -63 , 10),
  				conv_std_logic_vector( -75 , 10),
  				conv_std_logic_vector( -87 , 10),
  				conv_std_logic_vector(-100 , 10),
  				conv_std_logic_vector(-112 , 10),
  				conv_std_logic_vector(-124 , 10),
  				conv_std_logic_vector(-136 , 10),
  				conv_std_logic_vector(-148 , 10),
  				conv_std_logic_vector(-160 , 10),
  				conv_std_logic_vector(-172 , 10),
  				conv_std_logic_vector(-184 , 10),
  				conv_std_logic_vector(-196 , 10),
  				conv_std_logic_vector(-207 , 10),
  				conv_std_logic_vector(-218 , 10),
  				conv_std_logic_vector(-230 , 10),
  				conv_std_logic_vector(-241 , 10),
  				conv_std_logic_vector(-252 , 10),
  				conv_std_logic_vector(-263 , 10),
  				conv_std_logic_vector(-273 , 10),
  				conv_std_logic_vector(-284 , 10),
  				conv_std_logic_vector(-294 , 10),
  				conv_std_logic_vector(-304 , 10),
  				conv_std_logic_vector(-314 , 10),
  				conv_std_logic_vector(-324 , 10),
  				conv_std_logic_vector(-334 , 10),
  				conv_std_logic_vector(-343 , 10),
  				conv_std_logic_vector(-352 , 10),
  				conv_std_logic_vector(-361 , 10),
  				conv_std_logic_vector(-370 , 10),
  				conv_std_logic_vector(-379 , 10),
  				conv_std_logic_vector(-387 , 10),
  				conv_std_logic_vector(-395 , 10),
  				conv_std_logic_vector(-403 , 10),
  				conv_std_logic_vector(-410 , 10),
  				conv_std_logic_vector(-418 , 10),
  				conv_std_logic_vector(-425 , 10),
  				conv_std_logic_vector(-432 , 10),
  				conv_std_logic_vector(-438 , 10),
  				conv_std_logic_vector(-445 , 10),
  				conv_std_logic_vector(-451 , 10),
  				conv_std_logic_vector(-456 , 10),
  				conv_std_logic_vector(-462 , 10),
  				conv_std_logic_vector(-467 , 10),
  				conv_std_logic_vector(-472 , 10),
  				conv_std_logic_vector(-477 , 10),
  				conv_std_logic_vector(-481 , 10),
  				conv_std_logic_vector(-485 , 10),
  				conv_std_logic_vector(-489 , 10),
  				conv_std_logic_vector(-492 , 10),
  				conv_std_logic_vector(-496 , 10),
  				conv_std_logic_vector(-499 , 10),
  				conv_std_logic_vector(-501 , 10),
  				conv_std_logic_vector(-503 , 10),
  				conv_std_logic_vector(-505 , 10),
  				conv_std_logic_vector(-507 , 10),
  				conv_std_logic_vector(-509 , 10),
  				conv_std_logic_vector(-510 , 10),
  				conv_std_logic_vector(-510 , 10),
  				conv_std_logic_vector(-511 , 10),
  				conv_std_logic_vector(-511 , 10),
  				conv_std_logic_vector(-511 , 10),
  				conv_std_logic_vector(-510 , 10),
  				conv_std_logic_vector(-510 , 10),
  				conv_std_logic_vector(-509 , 10),
  				conv_std_logic_vector(-507 , 10),
  				conv_std_logic_vector(-505 , 10),
  				conv_std_logic_vector(-503 , 10),
  				conv_std_logic_vector(-501 , 10),
  				conv_std_logic_vector(-499 , 10),
  				conv_std_logic_vector(-496 , 10),
  				conv_std_logic_vector(-492 , 10),
  				conv_std_logic_vector(-489 , 10),
  				conv_std_logic_vector(-485 , 10),
  				conv_std_logic_vector(-481 , 10),
  				conv_std_logic_vector(-477 , 10),
  				conv_std_logic_vector(-472 , 10),
  				conv_std_logic_vector(-467 , 10),
  				conv_std_logic_vector(-462 , 10),
  				conv_std_logic_vector(-456 , 10),
  				conv_std_logic_vector(-451 , 10),
  				conv_std_logic_vector(-445 , 10),
  				conv_std_logic_vector(-438 , 10),
  				conv_std_logic_vector(-432 , 10),
  				conv_std_logic_vector(-425 , 10),
  				conv_std_logic_vector(-418 , 10),
  				conv_std_logic_vector(-410 , 10),
  				conv_std_logic_vector(-403 , 10),
  				conv_std_logic_vector(-395 , 10),
  				conv_std_logic_vector(-387 , 10),
  				conv_std_logic_vector(-379 , 10),
  				conv_std_logic_vector(-370 , 10),
  				conv_std_logic_vector(-361 , 10),
  				conv_std_logic_vector(-352 , 10),
  				conv_std_logic_vector(-343 , 10),
  				conv_std_logic_vector(-334 , 10),
  				conv_std_logic_vector(-324 , 10),
  				conv_std_logic_vector(-314 , 10),
  				conv_std_logic_vector(-304 , 10),
  				conv_std_logic_vector(-294 , 10),
  				conv_std_logic_vector(-284 , 10),
  				conv_std_logic_vector(-273 , 10),
  				conv_std_logic_vector(-263 , 10),
  				conv_std_logic_vector(-252 , 10),
  				conv_std_logic_vector(-241 , 10),
  				conv_std_logic_vector(-230 , 10),
  				conv_std_logic_vector(-218 , 10),
  				conv_std_logic_vector(-207 , 10),
  				conv_std_logic_vector(-196 , 10),
  				conv_std_logic_vector(-184 , 10),
  				conv_std_logic_vector(-172 , 10),
  				conv_std_logic_vector(-160 , 10),
  				conv_std_logic_vector(-148 , 10),
  				conv_std_logic_vector(-136 , 10),
  				conv_std_logic_vector(-124 , 10),
  				conv_std_logic_vector(-112 , 10),
  				conv_std_logic_vector(-100 , 10),
  				conv_std_logic_vector( -87 , 10),
  				conv_std_logic_vector( -75 , 10),
  				conv_std_logic_vector( -63 , 10),
  				conv_std_logic_vector( -50 , 10),
  				conv_std_logic_vector( -38 , 10),
  				conv_std_logic_vector( -25 , 10),
  				conv_std_logic_vector( -13 , 10),
  				conv_std_logic_vector(   0 , 10),
  				conv_std_logic_vector(  13 , 10),
  				conv_std_logic_vector(  25 , 10),
  				conv_std_logic_vector(  38 , 10),
  				conv_std_logic_vector(  50 , 10),
  				conv_std_logic_vector(  63 , 10),
  				conv_std_logic_vector(  75 , 10),
  				conv_std_logic_vector(  87 , 10),
  				conv_std_logic_vector( 100 , 10),
  				conv_std_logic_vector( 112 , 10),
  				conv_std_logic_vector( 124 , 10),
  				conv_std_logic_vector( 136 , 10),
  				conv_std_logic_vector( 148 , 10),
  				conv_std_logic_vector( 160 , 10),
  				conv_std_logic_vector( 172 , 10),
  				conv_std_logic_vector( 184 , 10),
  				conv_std_logic_vector( 196 , 10),
  				conv_std_logic_vector( 207 , 10),
  				conv_std_logic_vector( 218 , 10),
  				conv_std_logic_vector( 230 , 10),
  				conv_std_logic_vector( 241 , 10),
  				conv_std_logic_vector( 252 , 10),
  				conv_std_logic_vector( 263 , 10),
  				conv_std_logic_vector( 273 , 10),
  				conv_std_logic_vector( 284 , 10),
  				conv_std_logic_vector( 294 , 10),
  				conv_std_logic_vector( 304 , 10),
  				conv_std_logic_vector( 314 , 10),
  				conv_std_logic_vector( 324 , 10),
  				conv_std_logic_vector( 334 , 10),
  				conv_std_logic_vector( 343 , 10),
  				conv_std_logic_vector( 352 , 10),
  				conv_std_logic_vector( 361 , 10),
  				conv_std_logic_vector( 370 , 10),
  				conv_std_logic_vector( 379 , 10),
  				conv_std_logic_vector( 387 , 10),
  				conv_std_logic_vector( 395 , 10),
  				conv_std_logic_vector( 403 , 10),
  				conv_std_logic_vector( 410 , 10),
  				conv_std_logic_vector( 418 , 10),
  				conv_std_logic_vector( 425 , 10),
  				conv_std_logic_vector( 432 , 10),
  				conv_std_logic_vector( 438 , 10),
  				conv_std_logic_vector( 445 , 10),
  				conv_std_logic_vector( 451 , 10),
  				conv_std_logic_vector( 456 , 10),
  				conv_std_logic_vector( 462 , 10),
  				conv_std_logic_vector( 467 , 10),
  				conv_std_logic_vector( 472 , 10),
  				conv_std_logic_vector( 477 , 10),
  				conv_std_logic_vector( 481 , 10),
  				conv_std_logic_vector( 485 , 10),
  				conv_std_logic_vector( 489 , 10),
  				conv_std_logic_vector( 492 , 10),
  				conv_std_logic_vector( 496 , 10),
  				conv_std_logic_vector( 499 , 10),
  				conv_std_logic_vector( 501 , 10),
  				conv_std_logic_vector( 503 , 10),
  				conv_std_logic_vector( 505 , 10),
  				conv_std_logic_vector( 507 , 10),
  				conv_std_logic_vector( 509 , 10),
  				conv_std_logic_vector( 510 , 10),
  				conv_std_logic_vector( 510 , 10),
  				conv_std_logic_vector( 511 , 10));
  				

			constant SINROM_Table : ROM_TYPE := ROM_TYPE '( 

					conv_std_logic_vector(   0,10),
					conv_std_logic_vector(  13,10),
					conv_std_logic_vector(  25,10),
					conv_std_logic_vector(  38,10),
					conv_std_logic_vector(  50,10),
					conv_std_logic_vector(  63,10),
					conv_std_logic_vector(  75,10),
					conv_std_logic_vector(  87,10),
					conv_std_logic_vector( 100,10),
					conv_std_logic_vector( 112,10),
					conv_std_logic_vector( 124,10),
					conv_std_logic_vector( 136,10),
					conv_std_logic_vector( 148,10),
					conv_std_logic_vector( 160,10),
					conv_std_logic_vector( 172,10),
					conv_std_logic_vector( 184,10),
					conv_std_logic_vector( 196,10),
					conv_std_logic_vector( 207,10),
					conv_std_logic_vector( 218,10),
					conv_std_logic_vector( 230,10),
					conv_std_logic_vector( 241,10),
					conv_std_logic_vector( 252,10),
					conv_std_logic_vector( 263,10),
					conv_std_logic_vector( 273,10),
					conv_std_logic_vector( 284,10),
					conv_std_logic_vector( 294,10),
					conv_std_logic_vector( 304,10),
					conv_std_logic_vector( 314,10),
					conv_std_logic_vector( 324,10),
					conv_std_logic_vector( 334,10),
					conv_std_logic_vector( 343,10),
					conv_std_logic_vector( 352,10),
					conv_std_logic_vector( 361,10),
					conv_std_logic_vector( 370,10),
					conv_std_logic_vector( 379,10),
					conv_std_logic_vector( 387,10),
					conv_std_logic_vector( 395,10),
					conv_std_logic_vector( 403,10),
					conv_std_logic_vector( 410,10),
					conv_std_logic_vector( 418,10),
					conv_std_logic_vector( 425,10),
					conv_std_logic_vector( 432,10),
					conv_std_logic_vector( 438,10),
					conv_std_logic_vector( 445,10),
					conv_std_logic_vector( 451,10),
					conv_std_logic_vector( 456,10),
					conv_std_logic_vector( 462,10),
					conv_std_logic_vector( 467,10),
					conv_std_logic_vector( 472,10),
					conv_std_logic_vector( 477,10),
					conv_std_logic_vector( 481,10),
					conv_std_logic_vector( 485,10),
					conv_std_logic_vector( 489,10),
					conv_std_logic_vector( 492,10),
					conv_std_logic_vector( 496,10),
					conv_std_logic_vector( 499,10),
					conv_std_logic_vector( 501,10),
					conv_std_logic_vector( 503,10),
					conv_std_logic_vector( 505,10),
					conv_std_logic_vector( 507,10),
					conv_std_logic_vector( 509,10),
					conv_std_logic_vector( 510,10),
					conv_std_logic_vector( 510,10),
					conv_std_logic_vector( 511,10),
					conv_std_logic_vector( 511,10),
					conv_std_logic_vector( 511,10),
					conv_std_logic_vector( 510,10),
					conv_std_logic_vector( 510,10),
					conv_std_logic_vector( 509,10),
					conv_std_logic_vector( 507,10),
					conv_std_logic_vector( 505,10),
					conv_std_logic_vector( 503,10),
					conv_std_logic_vector( 501,10),
					conv_std_logic_vector( 499,10),
					conv_std_logic_vector( 496,10),
					conv_std_logic_vector( 492,10),
					conv_std_logic_vector( 489,10),
					conv_std_logic_vector( 485,10),
					conv_std_logic_vector( 481,10),
					conv_std_logic_vector( 477,10),
					conv_std_logic_vector( 472,10),
					conv_std_logic_vector( 467,10),
					conv_std_logic_vector( 462,10),
					conv_std_logic_vector( 456,10),
					conv_std_logic_vector( 451,10),
					conv_std_logic_vector( 445,10),
					conv_std_logic_vector( 438,10),
					conv_std_logic_vector( 432,10),
					conv_std_logic_vector( 425,10),
					conv_std_logic_vector( 418,10),
					conv_std_logic_vector( 410,10),
					conv_std_logic_vector( 403,10),
					conv_std_logic_vector( 395,10),
					conv_std_logic_vector( 387,10),
					conv_std_logic_vector( 379,10),
					conv_std_logic_vector( 370,10),
					conv_std_logic_vector( 361,10),
					conv_std_logic_vector( 352,10),
					conv_std_logic_vector( 343,10),
					conv_std_logic_vector( 334,10),
					conv_std_logic_vector( 324,10),
					conv_std_logic_vector( 314,10),
					conv_std_logic_vector( 304,10),
					conv_std_logic_vector( 294,10),
					conv_std_logic_vector( 284,10),
					conv_std_logic_vector( 273,10),
					conv_std_logic_vector( 263,10),
					conv_std_logic_vector( 252,10),
					conv_std_logic_vector( 241,10),
					conv_std_logic_vector( 230,10),
					conv_std_logic_vector( 218,10),
					conv_std_logic_vector( 207,10),
					conv_std_logic_vector( 196,10),
					conv_std_logic_vector( 184,10),
					conv_std_logic_vector( 172,10),
					conv_std_logic_vector( 160,10),
					conv_std_logic_vector( 148,10),
					conv_std_logic_vector( 136,10),
					conv_std_logic_vector( 124,10),
					conv_std_logic_vector( 112,10),
					conv_std_logic_vector( 100,10),
					conv_std_logic_vector(  87,10),
					conv_std_logic_vector(  75,10),
					conv_std_logic_vector(  63,10),
					conv_std_logic_vector(  50,10),
					conv_std_logic_vector(  38,10),
					conv_std_logic_vector(  25,10),
					conv_std_logic_vector(  13,10),
					conv_std_logic_vector(   0,10),
					conv_std_logic_vector( -13,10),
					conv_std_logic_vector( -25,10),
					conv_std_logic_vector( -38,10),
					conv_std_logic_vector( -50,10),
					conv_std_logic_vector( -63,10),
					conv_std_logic_vector( -75,10),
					conv_std_logic_vector( -87,10),
					conv_std_logic_vector(-100,10),
					conv_std_logic_vector(-112,10),
					conv_std_logic_vector(-124,10),
					conv_std_logic_vector(-136,10),
					conv_std_logic_vector(-148,10),
					conv_std_logic_vector(-160,10),
					conv_std_logic_vector(-172,10),
					conv_std_logic_vector(-184,10),
					conv_std_logic_vector(-196,10),
					conv_std_logic_vector(-207,10),
					conv_std_logic_vector(-218,10),
					conv_std_logic_vector(-230,10),
					conv_std_logic_vector(-241,10),
					conv_std_logic_vector(-252,10),
					conv_std_logic_vector(-263,10),
					conv_std_logic_vector(-273,10),
					conv_std_logic_vector(-284,10),
					conv_std_logic_vector(-294,10),
					conv_std_logic_vector(-304,10),
					conv_std_logic_vector(-314,10),
					conv_std_logic_vector(-324,10),
					conv_std_logic_vector(-334,10),
					conv_std_logic_vector(-343,10),
					conv_std_logic_vector(-352,10),
					conv_std_logic_vector(-361,10),
					conv_std_logic_vector(-370,10),
					conv_std_logic_vector(-379,10),
					conv_std_logic_vector(-387,10),
					conv_std_logic_vector(-395,10),
					conv_std_logic_vector(-403,10),
					conv_std_logic_vector(-410,10),
					conv_std_logic_vector(-418,10),
					conv_std_logic_vector(-425,10),
					conv_std_logic_vector(-432,10),
					conv_std_logic_vector(-438,10),
					conv_std_logic_vector(-445,10),
					conv_std_logic_vector(-451,10),
					conv_std_logic_vector(-456,10),
					conv_std_logic_vector(-462,10),
					conv_std_logic_vector(-467,10),
					conv_std_logic_vector(-472,10),
					conv_std_logic_vector(-477,10),
					conv_std_logic_vector(-481,10),
					conv_std_logic_vector(-485,10),
					conv_std_logic_vector(-489,10),
					conv_std_logic_vector(-492,10),
					conv_std_logic_vector(-496,10),
					conv_std_logic_vector(-499,10),
					conv_std_logic_vector(-501,10),
					conv_std_logic_vector(-503,10),
					conv_std_logic_vector(-505,10),
					conv_std_logic_vector(-507,10),
					conv_std_logic_vector(-509,10),
					conv_std_logic_vector(-510,10),
					conv_std_logic_vector(-510,10),
					conv_std_logic_vector(-511,10),
					conv_std_logic_vector(-511,10),
					conv_std_logic_vector(-511,10),
					conv_std_logic_vector(-510,10),
					conv_std_logic_vector(-510,10),
					conv_std_logic_vector(-509,10),
					conv_std_logic_vector(-507,10),
					conv_std_logic_vector(-505,10),
					conv_std_logic_vector(-503,10),
					conv_std_logic_vector(-501,10),
					conv_std_logic_vector(-499,10),
					conv_std_logic_vector(-496,10),
					conv_std_logic_vector(-492,10),
					conv_std_logic_vector(-489,10),
					conv_std_logic_vector(-485,10),
					conv_std_logic_vector(-481,10),
					conv_std_logic_vector(-477,10),
					conv_std_logic_vector(-472,10),
					conv_std_logic_vector(-467,10),
					conv_std_logic_vector(-462,10),
					conv_std_logic_vector(-456,10),
					conv_std_logic_vector(-451,10),
					conv_std_logic_vector(-445,10),
					conv_std_logic_vector(-438,10),
					conv_std_logic_vector(-432,10),
					conv_std_logic_vector(-425,10),
					conv_std_logic_vector(-418,10),
					conv_std_logic_vector(-410,10),
					conv_std_logic_vector(-403,10),
					conv_std_logic_vector(-395,10),
					conv_std_logic_vector(-387,10),
					conv_std_logic_vector(-379,10),
					conv_std_logic_vector(-370,10),
					conv_std_logic_vector(-361,10),
					conv_std_logic_vector(-352,10),
					conv_std_logic_vector(-343,10),
					conv_std_logic_vector(-334,10),
					conv_std_logic_vector(-324,10),
					conv_std_logic_vector(-314,10),
					conv_std_logic_vector(-304,10),
					conv_std_logic_vector(-294,10),
					conv_std_logic_vector(-284,10),
					conv_std_logic_vector(-273,10),
					conv_std_logic_vector(-263,10),
					conv_std_logic_vector(-252,10),
					conv_std_logic_vector(-241,10),
					conv_std_logic_vector(-230,10),
					conv_std_logic_vector(-218,10),
					conv_std_logic_vector(-207,10),
					conv_std_logic_vector(-196,10),
					conv_std_logic_vector(-184,10),
					conv_std_logic_vector(-172,10),
					conv_std_logic_vector(-160,10),
					conv_std_logic_vector(-148,10),
					conv_std_logic_vector(-136,10),
					conv_std_logic_vector(-124,10),
					conv_std_logic_vector(-112,10),
					conv_std_logic_vector(-100,10),
					conv_std_logic_vector( -87,10),
					conv_std_logic_vector( -75,10),
					conv_std_logic_vector( -63,10),
					conv_std_logic_vector( -50,10),
					conv_std_logic_vector( -38,10),
					conv_std_logic_vector( -25,10),
					conv_std_logic_vector( -13,10));
end NCO_ROM_package;


